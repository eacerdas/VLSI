module hello;
  initial
    begin
      $display("Test for the script");
      $finish;
    end
endmodule
	