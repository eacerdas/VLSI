interface intf_arbiter (input logic clk);

  	logic reset, req_0, req_1, gnt_0, gnt_1;
  
endinterface